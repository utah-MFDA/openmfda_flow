module thing((* type="flow" *)input [SIZE-1:0] beads_in,
               (* type="flow" *) output [SIZE-1:0]beads_out,
               (* type="flow" *)input [SIZE-1:0]cells_in,
               (* type="flow" *) output[SIZE-1:0] cells_out,
               (* type="flow" *) output [SIZE-1:0]collect,
               (* type="flow" *) input [SIZE-1:0]lysis_buffer_in,
               (* type="flow" *) output [SIZE-1:0]lysis_buffer_out,
               (* type="flow" *) input [SIZE-1:0]push_line,
               (* type="flow" *) output [SIZE-1:0]waste_out,
               (* type="ctrl" *) input collect_ctrl,
               lysis_in_ctrl, lysis_out_ctrl,
               push_ctrl,
               pump1, pump2, pump3,
               sep_ctrl,
               sieve_ctrl,
               waste_ctrl,
               beads_ctrl, cells_in_ctrl, cells_out_ctrl,
               (* type="flush" *) output collect_flush,
               lysis_in_flush, lysis_out_flush,
               push_flush,
               pump1_flush, pump2_flush, pump3_flush,
               sep_flush,
               sieve_flush,
               waste_flush,
               beads_flush, cells_in_flush, cells_out_flush);
parameter SIZE = 2;

mRNAiso_bank #(SIZE) bank(beads_in,
               beads_out,
               cells_in,
               cells_out,
               collect,
               lysis_buffer_in,
               lysis_buffer_out,
               push_line,
               waste_out,
               lysis_in_ctrl, lysis_out_ctrl,
               push_ctrl,
               pump1, pump2, pump3,
               sep_ctrl,
               sieve_ctrl,
               waste_ctrl,
               beads_ctrl, cells_in_ctrl, cells_out_ctrl,
               collect_flush,
               lysis_in_flush, lysis_out_flush,
               push_flush,
               pump1_flush, pump2_flush, pump3_flush,
               sep_flush,
               sieve_flush,
               waste_flush,
               beads_flush, cells_in_flush, cells_out_flush);
endmodule
