

YPressurePump soln1 1 2 pressure=100k
Ychannel soln1_channel 1 2 3 4 length=7.65m

YPressurePump soln2 5 6 pressure=100k chemConcentration=100m
Ychannel soln2_channel 5 6 7 8 length=3.24m


Ychannel output0 9 0 10 11 length=5.9m
Ychannel connect1 12 13 14 15 length=1.18m
Ychannel connect2 16 17 18 19 length=1.18m
Ychannel connect4 20 21 22 23 length=3.27m
Ychannel connect5 24 25 26 27 length=15.05m
Ychannel connect6 28 29 30 31 length=4.41m
Ychannel connect7 32 33 34 35 length=2.68m
Yserpentine_50px_0 serp1 3 12 4 14
Yserpentine_150px_0 serp2 13 16 15 18
Yserpentine_300px_0 serp3 7 20 8 22
Yserpentine_300px_0 serp4 21 24 23 26
Yserpentine_300px_0 serp5 25 28 27 30
Yserpentine_300px_0 serp6 29 36 31 37
Ydiffmix_25px_0 mix1 17 36 32 19 37 34
Yserpentine_300px_0 serp11 33 9 35 10


.tran 0.1m 1m
.print tran V(10)
.end


