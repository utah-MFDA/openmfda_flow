module demo (
    soln1,
    out
);

input   soln1;
output  out;
serpentine_150px_0   serp1   (.in_fluid(soln1), .out_fluid(out));
endmodule
