 
MACRO p_serpentine_2(L1.d, L2.d, turns.d)
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN p_serpentine_0 0 0 ;
  SIZE #L1 + 60# BY #L2*turns + 60# ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.5 29.5 30.5 30.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT #((turns+1)%2)*L1+29.5# #turns*L2+29.5# #((turns+1)%2)*L1+30.5# #turns*L2+30.5# ;
    END
  END out_fluid
  OBS
    LAYER met2 ;
      RECT 30 30 #L1+60# #L2*turns+60# ;
    LAYER met3 ;
      RECT 30 30 #L1+60# #L2*turns+60# ;
    LAYER met4 ;
      RECT 30 30 #L1+60# #L2*turns+60# ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END p_serpentine_0
