module thing((* type="flow" *) input [4:0] pad_prep_inlet,
             (* type="flow" *) input [SIZE-1:0] pad_ring_inlet,
             (* type="flow" *) output [1:0] pad_prep_outlet,
             (* type="flow" *) output [SIZE-1:0] pad_ring_outlet,
             (* type="flow" *) output [SIZE-1:0] pad_collect,
            (* type="flow" *) input pad_bead_in,
             (* type="ctrl" *) input [4:0] pad_ctrl_inlet,
             (* type="ctrl" *) input pad_ctrl_prep_inlet,
             pad_ctrl_v1, pad_ctrl_v2, pad_ctrl_sv1,
             pad_ctrl_stage_in,
             pad_ctrl_stage_out, pad_ctrl_sieve,
             pad_ctrl_collect,
             pad_ctrl_stage_inlet, pad_ctrl_stage_outlet, pad_ctrl_bead,
            pad_ctrl_prep_ringout,
             (* type="ctrl" *) input  [1:0] pad_ctrl_prep_outlet,
             (* type="ctrl" *) input [2:0] pad_pump,
             (* type="flush" *) output [4:0] pad_flush_inlet,
             (* type="flush" *) output pad_flush_prep_inlet,
             pad_flush_v1, pad_flush_v2, pad_flush_sv1,
             pad_flush_stage_in,
             pad_flush_stage_out, pad_flush_sieve,
             pad_flush_collect,
             pad_flush_stage_inlet, pad_flush_stage_outlet, pad_flush_bead,
            pad_flush_prep_ringout,
             (* type="flush" *) output [1:0] pad_flush_prep_outlet,
             (* type="flush" *) output [2:0] pad_flush_pump);
  parameter SIZE = 10;

      ChIP_pads #(SIZE) thingy(
      .pad_prep_inlet(pad_prep_inlet),
       .pad_ring_inlet(pad_ring_inlet),
       .pad_prep_outlet(pad_prep_outlet),
       .pad_ring_outlet(pad_ring_outlet),
       .pad_collect(pad_collect),
       .pad_bead_in(pad_bead_in),
       .pad_ctrl_inlet(pad_ctrl_inlet),
       .pad_ctrl_prep_inlet(pad_ctrl_prep_inlet),
       .pad_ctrl_v1(pad_ctrl_v1),
       .pad_ctrl_v2(pad_ctrl_v2),
       .pad_ctrl_sv1(pad_ctrl_sv1),
       .pad_ctrl_stage_in(pad_ctrl_stage_in),
       .pad_ctrl_stage_out(pad_ctrl_stage_out),
       .pad_ctrl_sieve(pad_ctrl_sieve),
       .pad_ctrl_collect(pad_ctrl_collect),
       .pad_ctrl_stage_inlet(pad_ctrl_stage_inlet),
       .pad_ctrl_stage_outlet(pad_ctrl_stage_outlet),
       .pad_ctrl_bead(pad_ctrl_bead),
       .pad_ctrl_prep_ringout(pad_ctrl_prep_ringout),
       .pad_ctrl_prep_outlet(pad_ctrl_prep_outlet),
       .pad_pump(pad_pump),
       .pad_flush_inlet(pad_flush_inlet),
       .pad_flush_prep_inlet(pad_flush_prep_inlet),
       .pad_flush_v1(pad_flush_v1),
       .pad_flush_v2(pad_flush_v2),
       .pad_flush_sv1(pad_flush_sv1),
       .pad_flush_stage_in(pad_flush_stage_in),
             .pad_flush_stage_out(pad_flush_stage_out),
       .pad_flush_sieve(pad_flush_sieve),
       .pad_flush_collect(pad_flush_collect),
       .pad_flush_stage_inlet(pad_flush_stage_inlet),
       .pad_flush_stage_outlet(pad_flush_stage_outlet),
       .pad_flush_bead(pad_flush_bead),
       .pad_flush_prep_ringout(pad_flush_prep_ringout),
       .pad_flush_prep_outlet(pad_flush_prep_outlet),
       .pad_flush_pump(pad_flush_pump));
endmodule
