../../../../pdks/h.r.3.3_pdk/distrib/1.0.0/h.r.3.3_merged.lef