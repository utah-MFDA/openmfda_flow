../pdk/distrib/0.0.2/h.r.3.3_pads.lef