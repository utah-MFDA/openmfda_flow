module top (
inout port_0_0,
inout port_0_1,
inout port_0_2,
inout port_0_3,
inout port_0_4,
inout port_0_5,
inout port_0_6,
inout port_0_7,
inout port_1_0,
inout port_1_1,
inout port_1_2,
inout port_1_3,
inout port_1_4,
inout port_1_5,
inout port_1_6,
inout port_1_7,
inout port_2_0,
inout port_2_1,
inout port_2_2,
inout port_2_3,
inout port_2_4,
inout port_2_5,
inout port_2_6,
inout port_2_7,
inout port_3_0,
inout port_3_1,
inout port_3_2,
inout port_3_3,
inout port_3_4,
inout port_3_5,
inout port_3_6,
inout port_3_7)

demo_50px device(.soln1(port_2_3),
            .soln2(port_2_5),
            .soln3(port_3_4),
            .out(port_3_3));

endmodule
