h.r.3.3_merged_0.0.2.lef