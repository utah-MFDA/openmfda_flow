../pdk/Components/p.m.8.k_merged.lef