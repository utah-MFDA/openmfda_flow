module thing((* type="flow" *)input [SIZE-1:0] beads_in,
               (* type="flow" *) output [SIZE-1:0]beads_out,
               (* type="flow" *)input [SIZE-1:0]cells_in,
               (* type="flow" *) output[SIZE-1:0] cells_out,
               (* type="flow" *) output [SIZE-1:0]collect,
               (* type="flow" *) input [SIZE-1:0]lysis_buffer_in,
               (* type="flow" *) output [SIZE-1:0]lysis_buffer_out,
               (* type="flow" *) input [SIZE-1:0]push_line,
               (* type="flow" *) output [SIZE-1:0]waste_out,
               (* type="ctrl" *) input collect_ctrl,
               lysis_in_ctrl, lysis_out_ctrl,
               push_ctrl,
               pump1, pump2, pump3,
               sep_ctrl,
               sieve_ctrl,
               waste_ctrl,
               beads_ctrl, cells_in_ctrl, cells_out_ctrl,
               (* type="flush" *) output collect_flush,
               lysis_in_flush, lysis_out_flush,
               push_flush,
               pump1_flush, pump2_flush, pump3_flush,
               sep_flush,
               sieve_flush,
               waste_flush,
               beads_flush, cells_in_flush, cells_out_flush);
parameter SIZE = 1;

mRNAiso_pads #(SIZE) bank(
.pad_beads_in(beads_in),
.pad_beads_out(beads_out),
.pad_cells_in(cells_in),
.pad_cells_out(cells_out),
.pad_collect(collect),
.pad_lysis_buffer_in(lysis_buffer_in),
.pad_lysis_buffer_out(lysis_buffer_out),
.pad_push_line(push_line),
.pad_waste_out(waste_out),
.pad_collect_ctrl(collect_ctrl),
.pad_lysis_in_ctrl(lysis_in_ctrl),
.pad_lysis_out_ctrl(lysis_out_ctrl),
.pad_push_ctrl(push_ctrl),
.pad_pump1(pump1),
.pad_pump2(pump2),
.pad_pump3(pump3),
.pad_sep_ctrl(sep_ctrl),
.pad_sieve_ctrl(sieve_ctrl),
.pad_waste_ctrl(waste_ctrl),
.pad_beads_ctrl(beads_ctrl),
.pad_cells_in_ctrl(cells_in_ctrl),
.pad_cells_out_ctrl(cells_out_ctrl),
.pad_collect_flush(collect_flush),
.pad_lysis_in_flush(lysis_in_flush),
.pad_lysis_out_flush(lysis_out_flush),
.pad_push_flush(push_flush),
.pad_pump1_flush(pump1_flush),
.pad_pump2_flush(pump2_flush),
.pad_pump3_flush(pump3_flush),
.pad_sep_flush(sep_flush),
.pad_sieve_flush(sieve_flush),
.pad_waste_flush(waste_flush),
.pad_beads_flush(beads_flush),
.pad_cells_in_flush(cells_in_flush),
.pad_cells_out_flush(cells_out_flush));
endmodule
