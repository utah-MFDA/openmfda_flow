../pdk/distrib/1.0.0/h.r.3.3_pads.lef